/*
a. The code is incorrect since it doesn't update the output whenever there's a 
	change in input